library verilog;
use verilog.vl_types.all;
entity congAND_vlg_check_tst is
    port(
        pin_name1       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end congAND_vlg_check_tst;
