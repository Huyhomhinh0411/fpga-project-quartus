library verilog;
use verilog.vl_types.all;
entity fullaader_vlg_vec_tst is
end fullaader_vlg_vec_tst;
