library verilog;
use verilog.vl_types.all;
entity congAND_vlg_vec_tst is
end congAND_vlg_vec_tst;
